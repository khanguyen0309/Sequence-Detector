//System Verilog testbench for 101 module
`timescale 1ns/1ps

module tb_101;
